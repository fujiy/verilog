module cpu ();

endmodule
